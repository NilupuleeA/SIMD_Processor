module addr_decoder (
    ports
);
    
endmodule
